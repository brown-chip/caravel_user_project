`default_nettype none

`timescale 1 ns / 1 ps

`include "uprj_netlists.v"
`include "caravel_netlists.v"

module cov_test_tb;
	

endmodule
`default_nettype wire
